`timescale 1ns / 1ps

module Mux_16X1_tb();
reg [15:0] I;
reg [3:0] S;
wire Y;

Mux_16X1 uut(.I(I), .S(S), .Y(Y));

initial begin
I = 16'b0000000000000000;  
     
        
I = 16'b0101011011010101; 
S = 4'b0000; 
#10;
S = 4'b0001; 
#10;
S = 4'b0010; 
#10;
S = 4'b0011; 
#10;
S = 4'b0100; 
#10;
S = 4'b0101; 
#10;
S = 4'b0110; 
#10;
S = 4'b0111; 
#10;
S = 4'b1000; 
#10;
S = 4'b1001; 
#10;
S = 4'b1010; 
#10;
S = 4'b1011; 
#10;
S = 4'b1100; 
#10;
S = 4'b1101; 
#10;
S = 4'b1110; 
#10;
S = 4'b1111; 
#10;
    
      
end

endmodule
