`timescale 1ns / 1ps

module Encoder_16X4_tb;

    reg [15:0] X;
    wire [3:0] Y;

    Encoder_16X4 uut (
        .X(X),
        .Y(Y)
    );

    initial begin
      
        X = 16'b0000000000000001; #10;
        X = 16'b0000000000000010; #10;
        X = 16'b0000000000000100; #10;
        X = 16'b0000000000001000; #10;
        X = 16'b0000000000010000; #10;
        X = 16'b0000000000100000; #10;
        X = 16'b0000000100000000; #10;
        X = 16'b0000001000000000; #10;
        X = 16'b0001000001000000; #10;
        X = 16'b0010000000000000; #10;
        X = 16'b0100000000100000; #10;
        X = 16'b1000010000000000; #10;
        X = 16'b1000010000100001; #10;
        X = 16'b0100000000011000; #10;
        X = 16'b0010000010000000; #10;
        X = 16'b1111000000000000; #10;
        X = 16'b0000111100000000; #10;
        X = 16'b0000000000110000; #10;
        X = 16'b0000000000001111; #10;
        X = 16'b1111111111111111; #10;
        X = 16'b0000000000000000; #10;

        $finish;
    end

endmodule
